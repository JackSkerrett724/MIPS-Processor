library ieee;
use ieee.std_logic_1164.all;
package globals is
constant BIT_WIDTH : integer := 8;
constant LOG_PORT_DEPTH : integer := 3;
end;

