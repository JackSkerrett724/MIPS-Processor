library ieee;
use ieee.std_logic_1164.all;
package globals is
constant N : INTEGER := 32;
constant M : INTEGER := 5;
end;

